* SPICE diode model for D1 in rct cellview
* .subckt DIODEM2 1 2
* D1 1 2 DIODEM2
.MODEL DIODEM2 D RS=1 CJO=0.1e-12
* .ends
